library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--library icai---impoertar libreria de paquete de constantes

package pkg_constant is
	constant R : integer := 
	constant I    "000"
	constant S    "
	constant B
	constant U
	constant J





--constant oor : std_logic_vector()